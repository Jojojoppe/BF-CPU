library IEEE;
use IEEE.STD_LOGIC_1164.all;
use work.all;

entity BF_CPU is
	port(
		CLK			: in std_logic;
		RST			: in std_logic;

		-- Debug output
		LED			: out std_logic_vector(7 downto 0)
	);
end entity;

architecture a of BF_CPU is
	-- Internal main signals
	signal nRST			: std_logic;		-- Inverted of RST (active high)
	signal sRST			: std_logic;		-- Software reset

	-- CPU lines
	signal CPU_D		: std_logic_vector(7 downto 0);
	signal CPU_A		: std_logic_vector(31 downto 0);

	-- RAM control lines
	signal RAM_wr		: std_logic;
	signal RAM_rd		: std_logic;

	-- Control lines registers
	signal AC_wr		: std_logic;	-- Accumulator
	signal AC_rd		: std_logic;
	signal IR_wr		: std_logic;	-- Instruction register
	signal IR_rd		: std_logic;

	-- Control lines pointer registers
	signal IP_wr		: std_logic;	-- Instruction pointer
	signal IP_rd		: std_logic;
	signal DP_wr		: std_logic;	-- Data pointer
	signal DP_rd		: std_logic;
	signal SP_wr		: std_logic;	-- Stack pointer
	signal SP_rd		: std_logic;

	-- Direct data lines
	signal AC_d			: std_logic_vector(7 downto 0);
	signal IR_d			: std_logic_vector(7 downto 0);
	signal IP_d			: std_logic_vector(31 downto 0);
	signal DP_d			: std_logic_vector(31 downto 0);
	signal SP_d			: std_logic_vector(31 downto 0);

	-- Arithmetic control lines
	signal DAR_inc		: std_logic;
	signal DAR_dec		: std_logic;
	signal AAR_inc		: std_logic;
	signal AAR_dec		: std_logic;
	signal AAR_adr		: std_logic_vector(31 downto 0);
	signal AAR_sel		: std_logic_vector(2 downto 0); -- Address arithmetic selector [IP, DP, SP]

	-- Data->Address bridge
	signal DAB_sel		: std_logic_vector(3 downto 0);
	signal DAB_en		: std_logic;
	signal DAB_d0		: std_logic_vector(7 downto 0);
	signal DAB_d1		: std_logic_vector(7 downto 0);
	signal DAB_d2		: std_logic_vector(7 downto 0);
	signal DAB_d3		: std_logic_vector(7 downto 0);

	-- Address->Data bridge
	signal ADB_sel		: std_logic_vector(3 downto 0);
	signal ADB_d0		: std_logic_vector(7 downto 0);
	signal ADB_d1		: std_logic_vector(7 downto 0);
	signal ADB_d2		: std_logic_vector(7 downto 0);
	signal ADB_d3		: std_logic_vector(7 downto 0);

	signal state		: integer;

begin

	-- Internal main signals
	nRST <= not(RST) or sRST;

	-- DEBUG LEDS
	LED <= CPU_D;

	-- Registers
	e_AC : entity REG8(a)			-- Accumulator
		port map(CLK, nRST, AC_rd, AC_wr, CPU_D, CPU_D, AC_d);
	e_IR : entity REG8(a)			-- Instruction register
		port map(CLK, nRST, IR_rd, IR_wr, CPU_D, CPU_D, IR_d);

	-- Data arithmetic (add/sub))
	e_DAR : entity INC8(a)
		port map(CLK, nRST, DAR_inc, DAR_dec, AC_d, CPU_d);

	-- Address arithmetic (add/sub)
	e_AARMux : entity MUX32_3(a)
		port map(CLK, nRST, AAR_sel, IP_d, DP_d, SP_d, AAR_adr);
	e_AAR : entity INC32(a)
		port map(CLK, nRST, AAR_inc, AAR_dec, AAR_adr, CPU_A);

	-- Pointer registers
	e_IP : entity REG32(a)			-- Instruction pointer
		port map(CLK, nRST, IP_rd, IP_wr, CPU_A, CPU_A, IP_d);
	e_DP : entity REG32(a)			-- Data pointer
		port map(CLK, nRST, DP_rd, DP_wr, CPU_A, CPU_A, DP_d);
	e_SP : entity REG32(a)			-- Data pointer
		port map(CLK, nRST, SP_rd, SP_wr, CPU_A, CPU_A, SP_d);

	-- Data->Address bridge
	e_DAB : entity DEMUX8_4(a)
		port map(CLK, nRST, DAB_sel, CPU_D, DAB_d0, DAB_d1, DAB_d2, DAB_d3);
	CPU_A <= DAB_d3 & DAB_d2 & DAB_d1 & DAB_d0 when (DAB_en = '1') else "ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ";

	-- Address->Data bridge
	e_ADB : entity MUX8_4(a)
		port map(CLK, nRST, ADB_sel, ADB_d0, ADB_d1, ADB_d2, ADB_d3, CPU_D);
	ADB_d0 <= CPU_A(7 downto 0);
	ADB_d1 <= CPU_A(15 downto 8);
	ADB_d2 <= CPU_A(23 downto 16);
	ADB_d3 <= CPU_A(31 downto 24);

	-- CONROL
	-- ------
	p_control : process(CLK, nRST)
	begin
		if nRST='1' then
			state <= 0;	-- Reset the CPU

		-- Control loop
		elsif rising_edge(CLK) then
			sRST		<= '0';

			AC_wr		<= '0';
			AC_rd		<= '0';
			IR_wr		<= '0';
			IR_rd		<= '0';
			IP_wr		<= '0';
			IP_rd		<= '0';
			DP_wr		<= '0';
			DP_rd		<= '0';
			SP_wr		<= '0';
			SP_rd		<= '0';

			DAR_inc		<= '0';
			DAR_dec		<= '0';
			AAR_inc		<= '0';
			AAR_dec		<= '0';
			AAR_sel		<= "000";

			DAB_sel		<= "0000";
			DAB_en		<= '0';

			ADB_sel		<= "0000";

			RAM_wr		<= '0';
			RAM_rd		<= '0';

			case state is

				-- Reset CPU
				when 0 =>
					state		<= 1;

				-- Fetch opcode from memory
				when 1 =>
					-- IR = RAM[IP]
					RAM_rd		<= '1';
					IR_wr		<= '1';
					IP_rd		<= '1';

					state		<= 2;

				-- Increase IP and decode opcode
				when 2 =>
					-- IP++
					IP_wr		<= '1';
					AAR_inc		<= '1';
					AAR_sel		<= "001";

					-- Decode opcode
					case IR_d(3 downto 0) is
						-- " " NOP
						when x"0" => state <= 1;
						-- ">" DP++
						when x"1" => state <= 3;
						-- "<" DP--
						when x"2" => state <= 4;
						-- "+" RAM[DP]++
						when x"3" => state <= 5;
						-- "-" RAM[DP] --
						when x"4" => state <= 7;
						-- "[" Conditional forward jump
						when x"5" => state <= 9;
						-- "]" Conditional backward jump
						when x"6" => state <= 14;
						-- Unknown -> RESET CPU
						when others =>
							sRST <= '0';
							state <= 0;
					end case;

				-- Increase DP
				when 3 =>
					-- DP++
					DP_wr		<= '1';
					AAR_sel		<= "010";
					AAR_inc		<= '1';
					state		<= 1;

				-- Decrease DP
				when 4 =>
					-- DP--
					DP_wr		<= '1';
					AAR_sel		<= "010";
					AAR_dec		<= '1';
					state		<= 2;

				-- Increase RAM[DP]
				when 5 =>
					-- AC = RAM[DP]
					RAM_rd		<= '1';
					AC_wr		<= '1';
					DP_rd		<= '1';
					state		<= 6;
				when 6 =>
					-- RAM[DP] = AC+1
					RAM_wr		<= '1';
					DAR_inc		<= '1';
					DP_rd		<= '1';
					state		<= 1;

				-- Decrease RAM[DP]
				when 7 =>
					-- AC = RAM[DP]
					RAM_rd		<= '1';
					AC_wr		<= '1';
					DP_rd		<= '1';
					state		<= 6;
				when 8 =>
					-- RAM[DP] = AC-1
					RAM_wr		<= '1';
					DAR_dec		<= '1';
					DP_rd		<= '1';
					state		<= 1;

				-- Conditional forward jump
				when 9 =>
					-- AC = RAM[DP]
					RAM_rd		<= '1';
					AC_wr		<= '1';
					DP_rd		<= '1';
					state		<= 10;
				when 10 =>
					-- Condition check
					if AC_d = x"00" then
						-- AC = IP[0]
						AC_wr		<= '1';
						ADB_sel		<= "0001";
						IP_rd		<= '1';
						state		<= 11;
					else
						-- AC = RAM[IP]
						RAM_rd		<= '1';
						IP_rd		<= '1';
						AC_wr		<= '1';
						state		<= 22;
				when 11 =>
					-- RAM[SP] = AC
					SP_rd		<= '1';
					RAM_wr		<= '1';
					AC_rd		<= '1';
					state		<= 12;
				when 12 =>
					-- SP--
					SP_wr		<= '1';
					AAR_sel		<= "100";
					AAR_dec		<= '1';
					state		<= 13;
				when 13 =>
					-- AC = IP[1]
					AC_wr		<= '1';
					ADB_sel		<= "0010";
					IP_rd		<= '1';
					state		<= 14;
				when 14 =>
					-- RAM[SP] = AC
					SP_rd		<= '1';
					RAM_wr		<= '1';
					AC_rd		<= '1';
					state		<= 15;
				when 15 =>
					-- SP--
					SP_wr		<= '1';
					AAR_sel		<= "100";
					AAR_dec		<= '1';
					state		<= 16;
				when 16 =>
					-- AC = IP[2]
					AC_wr		<= '1';
					ADB_sel		<= "0100";
					IP_rd		<= '1';
					state		<= 17;
				when 17 =>
					-- RAM[SP] = AC
					SP_rd		<= '1';
					RAM_wr		<= '1';
					AC_rd		<= '1';
					state		<= 18;
				when 18 =>
					-- SP--
					SP_wr		<= '1';
					AAR_sel		<= "100";
					AAR_dec		<= '1';
					state		<= 19;
				when 19 =>
					-- AC = IP[3]
					AC_wr		<= '1';
					ADB_sel		<= "1000";
					IP_rd		<= '1';
					state		<= 20;
				when 20 =>
					-- RAM[SP] = AC
					SP_rd		<= '1';
					RAM_wr		<= '1';
					AC_rd		<= '1';
					state		<= 21;
				when 21 =>
					-- SP--
					SP_wr		<= '1';
					AAR_sel		<= "100";
					AAR_dec		<= '1';
					state		<= 1;
				when 22 =>
					-- Check for ]
					if AC_d(3 downto 0) = x"6" then
						-- Execute ] (which will be NOP)
						state		<= 1;
					else
						-- IP++
						IP_wr		<= '1';
						AAR_sel		<= "001";
						AAR_inc		<= '1';
						state		<= 23;
				when 23 =>
					-- AC = RAM[IP]
					AC_wr		<= '1';
					RAM_rd		<= '1';
					IP_rd		<= '1';
					state		<= 22;

				-- Unknown state -> reset CPU
				when others =>
					sRST		<= '1';
					state		<= 0;
			end case;
		end if;
	end process;

end architecture;
